package yapp_pkj;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "./sv/yapp_packet.sv"
    `include "./sv/yapp_tx_monitor.sv"
    `include "./sv/yapp_tx_sequencer.sv"
    `include "./sv/yapp_tx_seqs.sv"
    `include "./sv/yapp_tx_driver.sv"
    `include "./sv/yapp_tx_agent.sv"
    `include "./sv/yap_env.sv"

endpackage: yapp_pkj